-- enmascarador.vhdl : Achivo VHDL generado automaticamente por el generador de c�digo RAILIB
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--entidad de enmascarador
entity enmascarador is
	generic(
		N_CVS : natural := 3;
		N_SEM : natural := 3;
		N_PAN : natural := 1;
		N_MDC : natural := 2;
		N_RUT : natural := 3
	);
	port(
		Clock : in std_logic;
		Reset : in std_logic;
		Modo : in std_logic_vector(N_RUT-1 downto 0);
		Ruta_in : in std_logic_vector(N_RUT-1 downto 0);
		Circuito_de_via : in std_logic_vector(N_CVS-1 downto 0);
		Semaforo_rojo_in : in std_logic_vector(N_SEM-1 downto 0);
		Semaforo_amarillo_in : in std_logic_vector(N_SEM-1 downto 0);
		Semaforo_verde_in : in std_logic_vector(N_SEM-1 downto 0);
		Barrera_alta_in : in std_logic_vector(N_PAN-1 downto 0);
		Barrera_baja_in : in std_logic_vector(N_PAN-1 downto 0);
		Maquina_normal_in : in std_logic_vector(N_MDC-1 downto 0);
		Maquina_reversa_in : in std_logic_vector(N_MDC-1 downto 0);
		Ocupacion : out std_logic_vector(N_CVS-1 downto 0);
		CV_int_Ruta_1 : out std_logic;
		CV_paralelo_Ruta_1 : out std_logic_vector(2-1 downto 0);
		CV_paralelo_temp_Ruta_1 : out std_logic_vector(3-1 downto 0);
		CV_despeje_Ruta_1 : out std_logic_vector(4-1 downto 0);
		CV_aprox_Ruta_1 : out std_logic_vector(5-1 downto 0);
		Estado_sub_ruta_Ruta_1 : out std_logic_vector(6-1 downto 0);
		Estado_ruta_cond_Ruta_1 : out std_logic_vector(7-1 downto 0);
		Estado_ruta_confl_Ruta_1 : out std_logic_vector(8-1 downto 0);
		Estado_SEM_sgte_Ruta_1 : out std_logic_vector(9-1 downto 0);
		Pos_MDC_ruta_Ruta_1 : out std_logic_vector(10-1 downto 0);
		Pos_MDC_aprox_Ruta_1 : out std_logic_vector(11-1 downto 0);
		Pos_MDC_despeje_Ruta_1 : out std_logic_vector(12-1 downto 0);
		Pos_MDC_solape_Ruta_1 : out std_logic_vector(13-1 downto 0);
		Bloq_MDC_ruta_Ruta_1 : out std_logic_vector(14-1 downto 0);
		Bloq_MDC_solape_Ruta_1 : out std_logic_vector(15-1 downto 0);
		Estado_PAN_Ruta_1 : out std_logic_vector(16-1 downto 0);
		Estado_CV_bloq_Ruta_1 : out std_logic;
		Estado_ruta_bloq_Ruta_1 : out std_logic_vector(18-1 downto 0);
		MDC_bloq_temp_solape_Ruta_1 : out std_logic_vector(19-1 downto 0);
		Estado_ruta_Ruta_1 : out std_logic_vector(20-1 downto 0);
		CV_alarma_total_Ruta_1 : out std_logic_vector(21-1 downto 0);
		CV_alarma_inmediata_Ruta_1 : out std_logic_vector(22-1 downto 0);
		PAN_bloq_temp_solape_Ruta_1 : out std_logic_vector(23-1 downto 0);
		CV_int_Ruta_2 : out std_logic;
		CV_paralelo_Ruta_2 : out std_logic_vector(2-1 downto 0);
		CV_paralelo_temp_Ruta_2 : out std_logic_vector(3-1 downto 0);
		CV_despeje_Ruta_2 : out std_logic_vector(4-1 downto 0);
		CV_aprox_Ruta_2 : out std_logic_vector(5-1 downto 0);
		Estado_sub_ruta_Ruta_2 : out std_logic_vector(6-1 downto 0);
		Estado_ruta_cond_Ruta_2 : out std_logic_vector(7-1 downto 0);
		Estado_ruta_confl_Ruta_2 : out std_logic_vector(8-1 downto 0);
		Estado_SEM_sgte_Ruta_2 : out std_logic_vector(9-1 downto 0);
		Pos_MDC_ruta_Ruta_2 : out std_logic_vector(10-1 downto 0);
		Pos_MDC_aprox_Ruta_2 : out std_logic_vector(11-1 downto 0);
		Pos_MDC_despeje_Ruta_2 : out std_logic_vector(12-1 downto 0);
		Pos_MDC_solape_Ruta_2 : out std_logic_vector(13-1 downto 0);
		Bloq_MDC_ruta_Ruta_2 : out std_logic_vector(14-1 downto 0);
		Bloq_MDC_solape_Ruta_2 : out std_logic_vector(15-1 downto 0);
		Estado_PAN_Ruta_2 : out std_logic_vector(16-1 downto 0);
		Estado_CV_bloq_Ruta_2 : out std_logic;
		Estado_ruta_bloq_Ruta_2 : out std_logic_vector(18-1 downto 0);
		MDC_bloq_temp_solape_Ruta_2 : out std_logic_vector(19-1 downto 0);
		Estado_ruta_Ruta_2 : out std_logic_vector(20-1 downto 0);
		CV_alarma_total_Ruta_2 : out std_logic_vector(21-1 downto 0);
		CV_alarma_inmediata_Ruta_2 : out std_logic_vector(22-1 downto 0);
		PAN_bloq_temp_solape_Ruta_2 : out std_logic_vector(23-1 downto 0);
		CV_int_Ruta_3 : out std_logic;
		CV_paralelo_Ruta_3 : out std_logic_vector(2-1 downto 0);
		CV_paralelo_temp_Ruta_3 : out std_logic_vector(3-1 downto 0);
		CV_despeje_Ruta_3 : out std_logic_vector(4-1 downto 0);
		CV_aprox_Ruta_3 : out std_logic_vector(5-1 downto 0);
		Estado_sub_ruta_Ruta_3 : out std_logic_vector(6-1 downto 0);
		Estado_ruta_cond_Ruta_3 : out std_logic_vector(7-1 downto 0);
		Estado_ruta_confl_Ruta_3 : out std_logic_vector(8-1 downto 0);
		Estado_SEM_sgte_Ruta_3 : out std_logic_vector(9-1 downto 0);
		Pos_MDC_ruta_Ruta_3 : out std_logic_vector(10-1 downto 0);
		Pos_MDC_aprox_Ruta_3 : out std_logic_vector(11-1 downto 0);
		Pos_MDC_despeje_Ruta_3 : out std_logic_vector(12-1 downto 0);
		Pos_MDC_solape_Ruta_3 : out std_logic_vector(13-1 downto 0);
		Bloq_MDC_ruta_Ruta_3 : out std_logic_vector(14-1 downto 0);
		Bloq_MDC_solape_Ruta_3 : out std_logic_vector(15-1 downto 0);
		Estado_PAN_Ruta_3 : out std_logic_vector(16-1 downto 0);
		Estado_CV_bloq_Ruta_3 : out std_logic;
		Estado_ruta_bloq_Ruta_3 : out std_logic_vector(18-1 downto 0);
		MDC_bloq_temp_solape_Ruta_3 : out std_logic_vector(19-1 downto 0);
		Estado_ruta_Ruta_3 : out std_logic_vector(20-1 downto 0);
		CV_alarma_total_Ruta_3 : out std_logic_vector(21-1 downto 0);
		CV_alarma_inmediata_Ruta_3 : out std_logic_vector(22-1 downto 0);
		PAN_bloq_temp_solape_Ruta_3 : out std_logic_vector(23-1 downto 0)
	);
end entity enmascarador;
-- Arquitectura del enmascarador : Descripcion del comportamiento
architecture enmascarador_ARQ of enmascarador is
	Signal Rojo_in_s,Amarillo_in_s,Verde_in_s,Rojo_out_s,Amarillo_out_s,Verde_out_s: std_logic_vector(N_SEM-1 downto 0);
	Signal Alto_in_s,Bajo_in_s,Alto_out_s,Bajo_out_s: std_logic_vector(N_PAN-1 downto 0);
	Signal Maquina_normal_in_s,Maquina_reversa_in_s,Maquina_normal_out_s,Maquina_reversa_out_s: std_logic_vector(N_MDC-1 downto 0);
	Signal Reset_sem_s,Reset_Pan_s: std_logic;
	begin
	process(Clock,Reset)
	begin
		if (Clock ='1' and Clock'Event) then
			if Reset = '1' then
				Estado_PAN_Ruta_1 <= (others => '0');
				PAN_bloq_temp_solape_Ruta_1 <= (others => '0');
				CV_alarma_inmediata_Ruta_1 <= (others => '0');
				CV_alarma_total_Ruta_1 <= (others => '0');
				CV_aprox_Ruta_1 <= (others => '0');
				CV_despeje_Ruta_1 <= (others => '0');
				CV_int_Ruta_1 <= '0';
				CV_paralelo_Ruta_1 <= (others => '0');
				CV_paralelo_temp_Ruta_1 <= (others => '0');
				MDC_bloq_temp_solape_Ruta_1 <= (others => '0');
				Pos_MDC_aprox_Ruta_1 <= (others => '0');
				Pos_MDC_despeje_Ruta_1 <= (others => '0');
				Pos_MDC_ruta_Ruta_1 <= (others => '0');
				Pos_MDC_solape_Ruta_1 <= (others => '0');
				Estado_ruta_Ruta_1 <= (others => '0');
				Estado_ruta_bloq_Ruta_1<= (others => '0');
				Estado_ruta_cond_Ruta_1<= (others => '0');
				Estado_ruta_confl_Ruta_1 <= (others => '0');
				Estado_sub_ruta_Ruta_1 <= (others => '0');
				Estado_SEM_sgte_Ruta_1 <= (others => '0');
				Estado_PAN_Ruta_2 <= (others => '0');
				PAN_bloq_temp_solape_Ruta_2 <= (others => '0');
				CV_alarma_inmediata_Ruta_2 <= (others => '0');
				CV_alarma_total_Ruta_2 <= (others => '0');
				CV_aprox_Ruta_2 <= (others => '0');
				CV_despeje_Ruta_2 <= (others => '0');
				CV_int_Ruta_2 <= '0';
				CV_paralelo_Ruta_2 <= (others => '0');
				CV_paralelo_temp_Ruta_2 <= (others => '0');
				MDC_bloq_temp_solape_Ruta_2 <= (others => '0');
				Pos_MDC_aprox_Ruta_2 <= (others => '0');
				Pos_MDC_despeje_Ruta_2 <= (others => '0');
				Pos_MDC_ruta_Ruta_2 <= (others => '0');
				Pos_MDC_solape_Ruta_2 <= (others => '0');
				Estado_ruta_Ruta_2 <= (others => '0');
				Estado_ruta_bloq_Ruta_2<= (others => '0');
				Estado_ruta_cond_Ruta_2<= (others => '0');
				Estado_ruta_confl_Ruta_2 <= (others => '0');
				Estado_sub_ruta_Ruta_2 <= (others => '0');
				Estado_SEM_sgte_Ruta_2 <= (others => '0');
				Estado_PAN_Ruta_3 <= (others => '0');
				PAN_bloq_temp_solape_Ruta_3 <= (others => '0');
				CV_alarma_inmediata_Ruta_3 <= (others => '0');
				CV_alarma_total_Ruta_3 <= (others => '0');
				CV_aprox_Ruta_3 <= (others => '0');
				CV_despeje_Ruta_3 <= (others => '0');
				CV_int_Ruta_3 <= '0';
				CV_paralelo_Ruta_3 <= (others => '0');
				CV_paralelo_temp_Ruta_3 <= (others => '0');
				MDC_bloq_temp_solape_Ruta_3 <= (others => '0');
				Pos_MDC_aprox_Ruta_3 <= (others => '0');
				Pos_MDC_despeje_Ruta_3 <= (others => '0');
				Pos_MDC_ruta_Ruta_3 <= (others => '0');
				Pos_MDC_solape_Ruta_3 <= (others => '0');
				Estado_ruta_Ruta_3 <= (others => '0');
				Estado_ruta_bloq_Ruta_3<= (others => '0');
				Estado_ruta_cond_Ruta_3<= (others => '0');
				Estado_ruta_confl_Ruta_3 <= (others => '0');
				Estado_sub_ruta_Ruta_3 <= (others => '0');
				Estado_SEM_sgte_Ruta_3 <= (others => '0');
			else
			Ocupacion(1) <= Ruta_in(1);
				Estado_PAN_Ruta_1(0) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(1) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(2) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(3) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(4) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(5) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(6) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(7) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(8) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(9) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(10) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(11) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(12) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(13) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_1(14) <= Barrera_alta_in(0);
				PAN_bloq_temp_solape_Ruta_1(0) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(1) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(2) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(3) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(4) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(5) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(6) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(7) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(8) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(9) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(10) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(11) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(12) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(13) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(14) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(15) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(16) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(17) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(18) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(19) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(20) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_1(21) <= Barrera_baja_in(0);
				CV_alarma_inmediata_Ruta_1(0) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_1(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(3) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(4) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_1(5) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(6) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(7) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_1(8) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(9) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(10) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(11) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(12) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_1(13) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(14) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_1(15) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(16) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(17) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(18) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_1(19) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_1(20) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_1(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(2) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_1(3) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(4) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(5) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_1(6) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(7) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_1(8) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(9) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(10) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(11) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(12) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_1(13) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_1(14) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(15) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(16) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(17) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_1(18) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_1(19) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_1(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_aprox_Ruta_1(1) <= Circuito_de_via(0);
				CV_aprox_Ruta_1(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_1(3) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_despeje_Ruta_1(0) <= Circuito_de_via(0);
				CV_despeje_Ruta_1(1) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_despeje_Ruta_1(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_int_Ruta_1 <= Circuito_de_via(0) or Circuito_de_via(1);
				Estado_CV_bloq_Ruta_1 <= Circuito_de_via(0) and Circuito_de_via(0);
				CV_paralelo_Ruta_1(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_paralelo_temp_Ruta_1(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_paralelo_temp_Ruta_1(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				MDC_bloq_temp_solape_Ruta_1(0) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(1) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(2) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(3) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(4) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(5) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(6) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(7) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(8) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(9) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(10) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(11) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(12) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(13) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(14) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(15) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(16) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_1(17) <= Maquina_reversa_in(0);
				Pos_MDC_aprox_Ruta_1(0) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(1) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(2) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(3) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(4) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(5) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(6) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(7) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(8) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_1(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(0) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(1) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(2) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(3) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(4) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(5) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(6) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(7) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(8) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_1(10) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(0) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(1) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(2) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(3) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(4) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(5) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(6) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(7) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_1(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(0) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(1) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(2) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(3) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(4) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(5) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(6) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(7) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(9) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(10) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_1(11) <= Maquina_normal_in(0);
				Estado_ruta_Ruta_1(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(1) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_1(2) <= Ruta_in(0);
				Estado_ruta_Ruta_1(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(4) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_1(5) <= Ruta_in(0);
				Estado_ruta_Ruta_1(6) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(7) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_1(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(9) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(10) <= Ruta_in(0);
				Estado_ruta_Ruta_1(11) <= Ruta_in(0);
				Estado_ruta_Ruta_1(12) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(13) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_1(14) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_1(15) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(16) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_1(17) <= Ruta_in(0);
				Estado_ruta_Ruta_1(18) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_1(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(5) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(6) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_1(7) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(9) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(10) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(11) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_1(12) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(13) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(14) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(15) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_1(16) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_1(0) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_1(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_1(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_1(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_1(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_1(5) <= Ruta_in(0);
				Estado_ruta_confl_Ruta_1(0) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(1) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(5) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_1(6) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_1(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_1(1) <= Ruta_in(0) or Ruta_in(2);
				Estado_sub_ruta_Ruta_1(2) <= Ruta_in(0) or Ruta_in(2);
				Estado_sub_ruta_Ruta_1(3) <= Ruta_in(0);
				Estado_sub_ruta_Ruta_1(4) <= Ruta_in(0) or Ruta_in(2);
				Bloq_MDC_ruta_Ruta_1(0) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(1) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(2) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(3) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(4) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(5) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(6) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(7) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(8) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(9) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(10) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_1(11) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_1(12) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_solape_Ruta_1(0) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(1) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(2) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(3) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(4) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(5) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(6) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_1(7) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(8) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(9) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(10) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_1(11) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_1(12) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_1(13) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Estado_SEM_sgte_Ruta_1(0) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1);
				Estado_SEM_sgte_Ruta_1(1) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_1(2) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_1(3) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1);
				Estado_SEM_sgte_Ruta_1(4) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1);
				Estado_SEM_sgte_Ruta_1(5) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_1(6) <= Semaforo_rojo_in(0);
				Estado_SEM_sgte_Ruta_1(7) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1);
				Estado_PAN_Ruta_2(0) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(1) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(2) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(3) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(4) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(5) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(6) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(7) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(8) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(9) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(10) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(11) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(12) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(13) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_2(14) <= Barrera_alta_in(0);
				PAN_bloq_temp_solape_Ruta_2(0) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(1) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(2) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(3) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(4) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(5) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(6) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(7) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(8) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(9) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(10) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(11) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(12) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(13) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(14) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(15) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(16) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(17) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(18) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(19) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(20) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_2(21) <= Barrera_baja_in(0);
				CV_alarma_inmediata_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_2(1) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(3) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(4) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_2(5) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(6) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(7) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(8) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_2(9) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(10) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(11) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_2(12) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(13) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(14) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(15) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_2(16) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(17) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(18) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(19) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_2(20) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_2(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(2) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_2(3) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(4) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(5) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(6) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_2(7) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(8) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_2(9) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(10) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(11) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(12) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(13) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(14) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(15) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(16) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(17) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(18) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_2(19) <= Circuito_de_via(0);
				CV_aprox_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_2(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_2(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_2(3) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_despeje_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_despeje_Ruta_2(1) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_despeje_Ruta_2(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_int_Ruta_2 <= Circuito_de_via(0) or Circuito_de_via(1);
				Estado_CV_bloq_Ruta_2 <= Circuito_de_via(0) and Circuito_de_via(0);
				CV_paralelo_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_paralelo_temp_Ruta_2(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_paralelo_temp_Ruta_2(1) <= Circuito_de_via(0);
				MDC_bloq_temp_solape_Ruta_2(0) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(1) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(2) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(3) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(4) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(5) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(6) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(7) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(8) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(9) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(10) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(11) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(12) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(13) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(14) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(15) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(16) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_2(17) <= Maquina_reversa_in(0);
				Pos_MDC_aprox_Ruta_2(0) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(1) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(2) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(3) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(4) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(5) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(6) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(7) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(8) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_2(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(0) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(1) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(2) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(3) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(4) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(5) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(6) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(7) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(8) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_2(10) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(0) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(1) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(2) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(3) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(4) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(5) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(6) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(7) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_2(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(0) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(1) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(2) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(3) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(4) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(5) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(6) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(7) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(9) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(10) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_2(11) <= Maquina_normal_in(0);
				Estado_ruta_Ruta_2(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_2(2) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_2(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(4) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_2(5) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_2(6) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(7) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_2(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(9) <= Ruta_in(0);
				Estado_ruta_Ruta_2(10) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_2(11) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(12) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_2(13) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(14) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(15) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(16) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(17) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_2(18) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_2(0) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(1) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(4) <= Ruta_in(0);
				Estado_ruta_bloq_Ruta_2(5) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(6) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_2(7) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(9) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(10) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(11) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(12) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(13) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_2(14) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_2(15) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_2(16) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_cond_Ruta_2(0) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_2(1) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_2(2) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_2(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_2(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_2(5) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_2(0) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_confl_Ruta_2(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_confl_Ruta_2(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_2(3) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_confl_Ruta_2(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_2(5) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_2(6) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_2(0) <= Ruta_in(0) or Ruta_in(1);
				Estado_sub_ruta_Ruta_2(1) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_2(2) <= Ruta_in(0) or Ruta_in(1);
				Estado_sub_ruta_Ruta_2(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_2(4) <= Ruta_in(0) or Ruta_in(1);
				Bloq_MDC_ruta_Ruta_2(0) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(1) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_2(2) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(3) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_2(4) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_2(5) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(6) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(7) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_2(8) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(9) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(10) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_2(11) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_2(12) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_solape_Ruta_2(0) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(1) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_2(2) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(3) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(4) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(5) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(6) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(7) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(8) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(9) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(10) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(11) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(12) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_2(13) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Estado_SEM_sgte_Ruta_2(0) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(1) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(2) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(3) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(4) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(5) <= Semaforo_rojo_in(0);
				Estado_SEM_sgte_Ruta_2(6) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_2(7) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_PAN_Ruta_3(0) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(1) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(2) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(3) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(4) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(5) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(6) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(7) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(8) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(9) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(10) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(11) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(12) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(13) <= Barrera_alta_in(0);
				Estado_PAN_Ruta_3(14) <= Barrera_alta_in(0);
				PAN_bloq_temp_solape_Ruta_3(0) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(1) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(2) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(3) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(4) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(5) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(6) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(7) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(8) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(9) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(10) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(11) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(12) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(13) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(14) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(15) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(16) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(17) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(18) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(19) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(20) <= Barrera_baja_in(0);
				PAN_bloq_temp_solape_Ruta_3(21) <= Barrera_baja_in(0);
				CV_alarma_inmediata_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_3(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(3) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(4) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_3(5) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(6) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_3(7) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(8) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(9) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(10) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_3(11) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_3(12) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(13) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(14) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(15) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_inmediata_Ruta_3(16) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(17) <= Circuito_de_via(0);
				CV_alarma_inmediata_Ruta_3(18) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(19) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_inmediata_Ruta_3(20) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(3) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(4) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(5) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(6) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(7) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(8) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(9) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(10) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(11) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_3(12) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(13) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(14) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_3(15) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_alarma_total_Ruta_3(16) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(17) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_alarma_total_Ruta_3(18) <= Circuito_de_via(0);
				CV_alarma_total_Ruta_3(19) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_3(1) <= Circuito_de_via(0);
				CV_aprox_Ruta_3(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_aprox_Ruta_3(3) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_despeje_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_despeje_Ruta_3(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_despeje_Ruta_3(2) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				CV_int_Ruta_3 <= Circuito_de_via(0) or Circuito_de_via(1);
				Estado_CV_bloq_Ruta_3 <= Circuito_de_via(0) and Circuito_de_via(0);
				CV_paralelo_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(1);
				CV_paralelo_temp_Ruta_3(0) <= Circuito_de_via(0) or Circuito_de_via(2);
				CV_paralelo_temp_Ruta_3(1) <= Circuito_de_via(0) or Circuito_de_via(1) or Circuito_de_via(2);
				MDC_bloq_temp_solape_Ruta_3(0) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(1) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(2) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(3) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(4) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(5) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(6) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(7) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(8) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(9) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(10) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(11) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(12) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(13) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(14) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(15) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(16) <= Maquina_reversa_in(0);
				MDC_bloq_temp_solape_Ruta_3(17) <= Maquina_reversa_in(0);
				Pos_MDC_aprox_Ruta_3(0) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(1) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(2) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(3) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(4) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(5) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(6) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(7) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(8) <= Maquina_normal_in(0);
				Pos_MDC_aprox_Ruta_3(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(0) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(1) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(2) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(3) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(4) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(5) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(6) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(7) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(8) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(9) <= Maquina_normal_in(0);
				Pos_MDC_despeje_Ruta_3(10) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(0) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(1) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(2) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(3) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(4) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(5) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(6) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(7) <= Maquina_normal_in(0);
				Pos_MDC_ruta_Ruta_3(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(0) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(1) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(2) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(3) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(4) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(5) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(6) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(7) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(8) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(9) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(10) <= Maquina_normal_in(0);
				Pos_MDC_solape_Ruta_3(11) <= Maquina_normal_in(0);
				Estado_ruta_Ruta_3(0) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_3(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_3(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(3) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_3(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(5) <= Ruta_in(0);
				Estado_ruta_Ruta_3(6) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(7) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_3(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(9) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_3(10) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_3(11) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(12) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_3(13) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(14) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_Ruta_3(15) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_Ruta_3(16) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(17) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_Ruta_3(18) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(1) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(4) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_3(5) <= Ruta_in(0);
				Estado_ruta_bloq_Ruta_3(6) <= Ruta_in(0);
				Estado_ruta_bloq_Ruta_3(7) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_3(8) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(9) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(10) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_3(11) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(12) <= Ruta_in(0);
				Estado_ruta_bloq_Ruta_3(13) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(14) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_bloq_Ruta_3(15) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_bloq_Ruta_3(16) <= Ruta_in(0);
				Estado_ruta_cond_Ruta_3(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_cond_Ruta_3(1) <= Ruta_in(0);
				Estado_ruta_cond_Ruta_3(2) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_cond_Ruta_3(3) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_cond_Ruta_3(4) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_cond_Ruta_3(5) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_3(0) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_3(1) <= Ruta_in(0) or Ruta_in(2);
				Estado_ruta_confl_Ruta_3(2) <= Ruta_in(0) or Ruta_in(1);
				Estado_ruta_confl_Ruta_3(3) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_3(4) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_ruta_confl_Ruta_3(5) <= Ruta_in(0);
				Estado_ruta_confl_Ruta_3(6) <= Ruta_in(0);
				Estado_sub_ruta_Ruta_3(0) <= Ruta_in(0) or Ruta_in(1);
				Estado_sub_ruta_Ruta_3(1) <= Ruta_in(0) or Ruta_in(1);
				Estado_sub_ruta_Ruta_3(2) <= Ruta_in(0) or Ruta_in(1) or Ruta_in(2);
				Estado_sub_ruta_Ruta_3(3) <= Ruta_in(0) or Ruta_in(1);
				Estado_sub_ruta_Ruta_3(4) <= Ruta_in(0) or Ruta_in(2);
				Bloq_MDC_ruta_Ruta_3(0) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(1) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_3(2) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_3(3) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(4) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(5) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_3(6) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_3(7) <= Maquina_reversa_in(0);
				Bloq_MDC_ruta_Ruta_3(8) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(9) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(10) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(11) <= Maquina_reversa_in(0) or Maquina_normal_in(1);
				Bloq_MDC_ruta_Ruta_3(12) <= Maquina_reversa_in(0);
				Bloq_MDC_solape_Ruta_3(0) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(1) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(2) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(3) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_3(4) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(5) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(6) <= Maquina_normal_in(0);
				Bloq_MDC_solape_Ruta_3(7) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(8) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(9) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(10) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(11) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(12) <= Maquina_normal_in(0) or Maquina_reversa_in(1);
				Bloq_MDC_solape_Ruta_3(13) <= Maquina_normal_in(0);
				Estado_SEM_sgte_Ruta_3(0) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_3(1) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_3(2) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_3(3) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1);
				Estado_SEM_sgte_Ruta_3(4) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_3(5) <= Semaforo_rojo_in(0);
				Estado_SEM_sgte_Ruta_3(6) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
				Estado_SEM_sgte_Ruta_3(7) <= Semaforo_rojo_in(0) or Semaforo_rojo_in(1) or Semaforo_amarillo_in(1) or Semaforo_verde_in(1) or Semaforo_rojo_in(2) or Semaforo_amarillo_in(2) or Semaforo_verde_in(2);
			end if;
		end if;
	end process;
end architecture enmascarador_ARQ;
