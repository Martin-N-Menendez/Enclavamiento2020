library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


-- AGREGAR salida que mate paquete_ok;

entity registro is
	port(
		clk_i: in std_logic;
        rst_i: in std_logic;
        procesar : in std_logic;
        procesado : out std_logic;
        paquete_i: in std_logic_vector(15-1 downto 0);
        w_data: out std_logic_vector(8-1 downto 0);
        wr_uart : out std_logic  -- "char_disp"
	);
    end entity;

architecture Behavioral of registro is
    
    type estados_t is (REINICIO,CICLO_1,CICLO_2);
    signal estado, estado_siguiente : estados_t;
  

    --signal paquete_aux: std_logic_vector(15-1 downto 0);
    signal mux_out_s : std_logic;
    signal ena_s : std_logic;
    signal rst_s : std_logic;  
    signal mux_s : std_logic_vector(4-1 downto 0);

   
begin    
   --<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<
    contador : process(clk_i)
    begin
        if (clk_i = '1' and clk_i'event) then
            if rst_i = '1' then
                mux_s <= "0000";
            elsif (ena_s = '1') then        
               if (mux_s = "1111") then
                   mux_s <= "0000";
               else
                   mux_s <= std_logic_vector(to_unsigned(to_integer(unsigned(mux_s)) + 1 , 4));         
               end if;
            end if; 
        end if;
    end process;
    
    multiplexor : process(paquete_i,mux_s)
    begin
        case mux_s is
            when "0000" => mux_out_s <= paquete_i(0);
            when "0001" => mux_out_s <= paquete_i(1);
            when "0010" => mux_out_s <= paquete_i(2);
            when "0011" => mux_out_s <= paquete_i(3);
            when "0100" => mux_out_s <= paquete_i(4);
            when "0101" => mux_out_s <= paquete_i(5);
            when "0110" => mux_out_s <= paquete_i(6);
            when "0111" => mux_out_s <= paquete_i(7);
            when "1000" => mux_out_s <= paquete_i(8);
            when "1001" => mux_out_s <= paquete_i(9);
            when "1010" => mux_out_s <= paquete_i(10);
            when "1011" => mux_out_s <= paquete_i(11);
            when "1100" => mux_out_s <= paquete_i(12);
            when "1101" => mux_out_s <= paquete_i(13);
            when "1110" => mux_out_s <= paquete_i(14);
            when others => mux_out_s <= '0';
        end case;
        
    end process;
    
--    bit_to_ascii : process(clk_i)
--    begin
--        if (clk_i = '1' and clk_i'event) then
--            if rst_i = '1' then
--                w_data <= (others => '0');
--            else                     
               w_data <= "00110001" when mux_out_s = '1' else "00110000";
--            end if; 
--    end process;
    
    FSM_reset : process(clk_i)
    begin
        if (clk_i = '1' and clk_i'event) then
            if rst_i = '1' then
                estado <= reinicio;          
            else          
               estado <= estado_siguiente;
            end if; 
        end if;
    end process;
    
    FSM : process(procesar,estado,mux_s)
    begin
        estado_siguiente <= estado;
        
        case estado is
            when REINICIO =>
                wr_uart <= '0';
                rst_s <= '1';
                ena_s <= '0';
                procesado <= '0';
                
                if procesar = '1' then
                    estado_siguiente <= CICLO_1;
                end if;
                
            when CICLO_1 =>
                wr_uart <= '0';
                rst_s <= '0';
                ena_s <= '0';
                --procesado <= '0';
                
                estado_siguiente <= CICLO_2;
                
            when CICLO_2 =>
                wr_uart <= '1';
                rst_s <= '0';
                ena_s <= '1';              
                procesado <= '0';
                
                if mux_s = "1110" then
                    procesado <= '1';
                    estado_siguiente <= REINICIO;           
                else
                    estado_siguiente <= CICLO_1;

                end if;
            when others => null;
        end case;
    end process;
        
end Behavioral;
