library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity conector_test is
	port(
		clk_i: in std_logic;
        rst_i: in std_logic;
        switch : in std_logic;
        leds : out std_logic_vector(2-1 downto 0);
        wr_uart_3 : out std_logic;
        N_1 : in integer;
        N_2 : in integer;
        r_disponible : in std_logic;
        w_data_1: in std_logic_vector(8-1 downto 0);
        w_data_2: in std_logic_vector(8-1 downto 0);
        w_data_3: out std_logic_vector(8-1 downto 0)
	);
    end entity;

architecture Behavioral of conector_test is
  
  signal disp_aux_1 : std_logic_vector(8-1 downto 0);
  signal disp_aux_2 : std_logic_vector(8-1 downto 0);
  signal disp_aux_3 : std_logic_vector(8-1 downto 0);
  signal disp_aux_4 : std_logic_vector(8-1 downto 0);
        
begin
     
    process(clk_i)
    variable contador: integer := 0;
    variable N_total : integer := 0;
    begin
        if (clk_i = '1' and clk_i'event) then
            if rst_i = '1' then
                N_total := 0; 
                contador := 0; 
            else 
                if switch = '1' then                 
                    
                    disp_aux_2 <= w_data_2;
                    
                    w_data_3 <= disp_aux_2;
                                 
                    wr_uart_3 <= r_disponible;
            
                    
                    --leds <= "10";
                else   
 
       
                    disp_aux_1 <= w_data_1;
                    
                    w_data_3 <= disp_aux_1;
                                 
                    wr_uart_3 <= r_disponible;
                        
     
                                       
      
                    --leds <= "01";
                end if;
            end if;
        end if;
    end process;  
    
        
end Behavioral;